module FFT#(parameter WIDTH=32,SIZE=32)(
	input []
);
