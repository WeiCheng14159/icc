module avg(din, reset, clk, ready, dout);
input reset, clk;
input [15:0] din;
output reg ready; 
output reg [15:0] dout;

// ==========================================
//  Enter your design below
// ==========================================



endmodule
